library verilog;
use verilog.vl_types.all;
entity sdram_ctrl_top_tst is
end sdram_ctrl_top_tst;
